module inst_mem(input [15:0] PC ,input en, output [15:0] instr);

reg [15:0] rom [65535:0];  
//integer i;
//

////////////////////////////////////////////////
//////////Testing Branch Predictor//////////////
////////////////////////////////////////////////
//initial begin
//rom[0] = 16'b0011011000001000;       //LLI 0011 011 000 001 000   r(3) = 8
//rom[1] = 16'b0011101000001000;       //LLI 0011 101 000 010 000   r(5) = 8
//rom[2] = 16'b0011100000001000;       //LLI 0011 100 000 010 000   r(4) = 8
//rom[3] = 16'b1000100011000011;        //BEQ 1000 101 011 010010  PC = 18*2
//rom[4] = 16'b0011101000001001;        //LLI 0011 101 000 010 000   r(5) = 9
//rom[5] = 16'b0011101000001011;        //LLI 0011 101 000 010 000   r(5) = 11
//rom[6] = 16'b0011101000001100;        //LLI 0011 101 000 010 000   r(5) = 12
//rom[7] = 16'b0011101000001100;        //LLI 0011 101 000 010 000   r(5) = 12
//rom[8] = 16'b0011101000001100;        //LLI 0011 101 000 010 000   r(5) = 12
//rom[9] = 16'b1011010111111000;       // JAL 1011 010 000000010    
////rom[7] = 16'b1000100011000011;        //using same brach instruction
////rom[10] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 11


//end

initial begin
rom[0] = 16'b0011011000001000;       //LLI 0011 011 000 001 000   r(3) = 8
rom[1] = 16'b0011101000001000;       //LLI 0011 101 000 010 000   r(5) = 8
rom[2] = 16'b0011100000001000;       //LLI 0011 100 000 010 000   r(4) = 8 //hump comes here
rom[3] = 16'b1000100011000010;        //BEQ 1000 101 011 010010  
rom[4] = 16'b0011101000001001;        //LLI 0011 101 000 010 000   r(5) = 9
rom[5] = 16'b0011101000001011;        //LLI 0011 101 000 010 000   r(5) = 11 //branch ccmes here
rom[6] = 16'b1000100011000011;        //BEQ 1000 101 011 010010  
rom[7] = 16'b0011101000001101;        //LLI 0011 101 000 010 000   r(5) = 12
rom[8] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 15
rom[9] = 16'b0011101000001101;        //LLI 0011 101 000 010 000   r(5) = 13 //brach comes here
rom[10]= 16'b1000100011000011;        //BEQ 1000 101 011 010010     
rom[11] = 16'b0011101000001100;        //LLI 0011 101 000 010 000   r(5) = 12
rom[12] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 15
rom[13] = 16'b0011101000000001;       //LLI 0011 101 000 010 000   r(5) = 1 //branch comes hers
rom[14] = 16'b0011101000001101;        //LLI 0011 101 000 010 000   r(5) = 13
rom[15] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 15
rom[16] = 16'b0011101000001101;        //LLI 0011 101 000 010 000   r(5) = 13
rom[17] = 16'b1011010111110001;       // JAL 1011 010 000000010
end
//initial begin 
////rom[0] = 16'b0011011000001000;       //LLI 0011 011 000 001 000   r(3) = 8
////rom[1] = 16'b0011101000001001;       //LLI 0011 101 000 010 000   r(5) = 9
////rom[2] = 16'b0011100000001010;       //LLI 0011 100 000 010 000   r(4) = 10
////rom[3] = 16'b0000011101110000;       // ADD 0000 011 101 110 000  r(6) = r(3) + r(5)
////rom[4] = 16'b0110101011011000;       //LM 0110 101 011011000 
////rom[5] = 16'b0000011101110000;       // ADD 0000 011 101 110 000  r(6) = r(3) + r(5)
//// to test branch and jump
//rom[0] = 16'b0011011000001000;       //LLI 0011 011 000 001 000   r(3) = 8
//rom[1] = 16'b0011101000001000;       //LLI 0011 101 000 010 000   r(5) = 8
//rom[3] = 16'b0011100000001000;       //LLI 0011 100 000 010 000   r(4) = 8
//rom[4] = 16'b1000100011000011;        //BEQ 1000 100 011 010010  PC = 18*2 //jump comes here
//rom[5] = 16'b0011101000001001;        //LLI 0011 101 000 010 000   r(5) = 9
//rom[6] = 16'b0011101000001011;        //LLI 0011 101 000 010 000   r(5) = 11
//rom[7] = 16'b0011101000001100;        //LLI 0011 101 000 010 000   r(5) = 12 //branch comes here
//rom[8] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 15
//rom[9] = 16'b0011101000001101;        //LLI 0011 101 000 010 000   r(5) = 13
////rom[10] = 16'b1011010111111010;       // JAL 1011 010 000000010    //jumps goes to 4 
//rom[10] = 16'b1011010111110110;       // JAL 1011 010 000000010    //jumps goes to 3 
////rom[7] = 16'b1000100011000011;        //using same brach instruction
////rom[10] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 11
//end


//initial begin
//initial begin
////LM and SM testing
//rom[0] = 16'b0011011000001000;       //LLI 0011 011 000 001 000   r(3) = 8
//rom[1] = 16'b0011101000001001;       //LLI 0011 101 000 001 001   r(5) = 9
//rom[2] = 16'b0011100000001000;       //LLI 0011 100 000 001 010   r(4) = 10
//rom[3] = 16'b0000011101110000;       // ADD 0000 011 101 110 000  r(6) = r(3) + r(5)
//rom[4] = 16'b0110101011011000;       //LM 0110 101 011011000 Load into r(7), r(6), r(4) and r(3)
//rom[5] = 16'b0000011101110000;       // ADD 0000 011 101 110 000  r(6) = r(3) + r(5)
//rom[6] = 16'b0111110001111000;       // SM 0111 110 001111000 store from r(6),r(5), r(4) and r(3)

////// to test branch and jump
////rom[3] = 16'b1000100011000011;        //BEQ 1000 100 011 010010  PC = 18*2
////rom[4] = 16'b0011101000001001;        //LLI 0011 101 000 010 000   r(5) = 9
////rom[5] = 16'b0011101000001011;        //LLI 0011 101 000 010 000   r(5) = 11
////rom[6] = 16'b0011101000001100;        //LLI 0011 101 000 010 000   r(5) = 12
////rom[7] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 15
////rom[8] = 16'b0011101000001101;        //LLI 0011 101 000 010 000   r(5) = 13
////rom[9] = 16'b1011010111111010;       // JAL 1011 010 000000010    
////rom[10] = 16'b1000100011000011;        //using same brach instruction
////rom[11] = 16'b0011101000001111;        //LLI 0011 101 000 010 000   r(5) = 11


//end
//////////////////////////////////////////////////////
///////////////Universal Code To Verify///////////////
//////////////////////////////////////////////////////
//initial begin
//rom[0] = 16'b0011011000001000;       //LLI 0011 011 000 001 000   r(3) = 8
//rom[1] = 16'b0011100000001000;       //LLI 0011 100 000 001 000   r(4) = 8
//rom[2] = 16'b0000011100110000;       //ADD 0000 011 101 110 000  r(6) = r(3) + r(4)
//rom[3] = 16'b1000100011000010;       //BEQ 1000 100 011 000011  target PC = 3 + 2
//rom[4] = 16'b0011101000001001;       //LLI 0011 101 000 001 001   r(5) = 9
//rom[5] = 16'b0011101000001000;       //LLI 0011 101 000 001 000   r(5) = 8 //comes here if branch at rom[3] is taken
//rom[6] = 16'b0110101011011000;       //LM 0110 101 011011000
//rom[7] = 16'b0000011101110000;       //ADD 0000 011 101 110 000  r(6) = r(3) + r(5)
//rom[8] = 16'b0111110001111000;       // SM 0111 110 001111000
//rom[9] = 16'b1011010111111001;       // JAL 1011 010 000000010

//end






assign instr = en ? rom[PC]:16'd0;
endmodule